`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:31:00 05/17/2012 
// Design Name: 
// Module Name:    shadow_capture_v2 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module shadow_capture_v2(
    input clk,
    input rst,
    input c_en,
    input d_clk,
    input [0:0] d_in,
    output [0:0] d_out,
    output d_ready
    );


endmodule
